`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Name: Loc Nguyen
// Course: ELC 5312
// Assignment: CR1
// Date: 9/11/2025
//////////////////////////////////////////////////////////////////////////////////


module top(
// port declaration 
    input  logic        clk_100mhz,   // Basys3 has clock of 100 MHz
    input  logic        rst_n,  // mapped to U18
    
    input  logic        en,           // enable circulation (1 = run, 0 = pause)
    input  logic        cw,           // 1 = clockwise, 0 = counter-clockwise
    output logic [6:0]  seg,          // segments a..g (active LOW)
    output logic        dp,           // decimal point (active LOW)
    output logic [3:0]  an            // anode enables (active LOW)
);
 logic rst_n_int;
    assign rst_n_int = ~rst_n;

    // ----------------------------------------------------------------
    // Timing parameters 
    // ----------------------------------------------------------------
    // ~1 kHz rate for digit scan. Calculation is 100_000_000 / 1khz = 100_000 is our division
    localparam int SCAN_DIV = 100_000;     // gives ~1 kHz digit refresh about 250 hz per digit

    // step rate 1 hz or every 1 second. Calculation 100_000_000/1hz = 100_000_000
    localparam int STEP_DIV = 100_000_000; // 1 step per second
    // ----------------------------------------------------------------
    // Clock dividers: scan tick for digit multiplexing, step tick for motion
    // ----------------------------------------------------------------
    logic [$clog2(SCAN_DIV)-1:0] scan_cnt = '0;
    logic                         scan_tick;
  
    always_ff @(posedge clk_100mhz or negedge rst_n_int) begin
        if (!rst_n_int) begin
            scan_cnt  <= '0;
            scan_tick <= 1'b0;
        end else begin
            if (scan_cnt == SCAN_DIV-1) begin
                scan_cnt  <= '0;
                scan_tick <= 1'b1;
            end else begin
                scan_cnt  <= scan_cnt + 1;
                scan_tick <= 1'b0;
            end
        end
    end

    logic [$clog2(STEP_DIV)-1:0] step_cnt = '0;
    logic                         step_tick;
    

    always_ff @(posedge clk_100mhz or negedge rst_n_int) begin
        if (!rst_n_int) begin
            step_cnt  <= '0;
            step_tick <= 1'b0;
        end else begin
            if (step_cnt == STEP_DIV-1) begin
                step_cnt  <= '0;
                step_tick <= 1'b1;
            end else begin
                step_cnt  <= step_cnt + 1;
                step_tick <= 1'b0;
            end
        end
    end

    // ----------------------------------------------------------------
    // 8-position state machine 
    // Sequence (clockwise):
    //   0: D0 top   -> 1: D1 top -> 2: D2 top -> 3: D3 top
    //   4: D3 bottom-> 5: D2 bottom -> 6: D1 bottom -> 7: D0 bottom -> back to 0
    // Counterclockwise is reverse order.
    // ----------------------------------------------------------------
    logic [2:0] state = 3'd0;

    function automatic [2:0] next_state(input [2:0] s, input logic cw_f);
        if (cw_f) begin
            next_state = (s == 3'd7) ? 3'd0 : s + 3'd1;
        end else begin
            next_state = (s == 3'd0) ? 3'd7 : s - 3'd1;
        end
    endfunction

    always_ff @(posedge clk_100mhz or negedge rst_n_int) begin
        if (!rst_n_int) begin
            state <= 3'd0;
        end else if (step_tick && en) begin
            state <= next_state(state, cw);
        end
    end

    // ----------------------------------------------------------------
    // Digit scanner 
    // ----------------------------------------------------------------
    logic [1:0] cur_digit = 2'd0; //2 bits counter values 0-3 for 4 digits
    always_ff @(posedge clk_100mhz or negedge rst_n_int) begin
        if (!rst_n_int) begin //reset behavior 
            cur_digit <= 2'd0; // if !rst_n then cur_digit = 0 start right most digit
        end else if (scan_tick) begin //slow clock enable pulse generated by dividing 100Mhz down to 1Khz
            cur_digit <= cur_digit + 2'd1; // for ea scan_tick = 1, cur_digit increment by 1 it does this from 0 to 3 then back to 0.
        end
    end

    // Active-LOW anode 
    always_comb begin
        an = 4'b1111;
        unique case (cur_digit)
            2'd0: an = 4'b1110; // enable digit 0 (rightmost on Basys3�s silkscreen)
            2'd1: an = 4'b1101; // digit 1
            2'd2: an = 4'b1011; // digit 2
            2'd3: an = 4'b0111; // digit 3 (leftmost)
        endcase
    end

    // ----------------------------------------------------------------
    // Segment patterns (active-LOW)
    // seg[6:0] = {a,b,c,d,e,f,g} with 0=ON
    // ----------------------------------------------------------------
    localparam logic [6:0] SEG_TOP_SQ    = 7'b0011100; //a = on, b = on, f = on, g = on
    localparam logic [6:0] SEG_BOT_SQ    = 7'b0100011; // g = on, c = on, d = on, e = on

    // bit6 g, bit5 b, bit4 c, bit3 d, bit2 e, bit1 f, bit0 a

 
    function automatic logic [6:0] square_for(input [2:0] s, input [1:0] digit);
       
        square_for = 7'b111_1111; //1 means anode is off

        // Map states to (digit, top/bottom)
        // 0: d0 top, 1: d1 top, 2: d2 top, 3: d3 top,
        // 4: d3 bot, 5: d2 bot, 6: d1 bot, 7: d0 bot
        unique case (s)
            3'd0: if (digit == 2'd0) square_for = SEG_TOP_SQ;
            3'd1: if (digit == 2'd1) square_for = SEG_TOP_SQ;
            3'd2: if (digit == 2'd2) square_for = SEG_TOP_SQ;
            3'd3: if (digit == 2'd3) square_for = SEG_TOP_SQ;
            3'd4: if (digit == 2'd3) square_for = SEG_BOT_SQ;
            3'd5: if (digit == 2'd2) square_for = SEG_BOT_SQ;
            3'd6: if (digit == 2'd1) square_for = SEG_BOT_SQ;
            3'd7: if (digit == 2'd0) square_for = SEG_BOT_SQ;
            default: /* keep blank */;
        endcase
    endfunction

    // Drive segments for the currently digit
    always_comb begin
        seg = square_for(state, cur_digit);
        dp  = 1'b1; // means always OFF
    end

endmodule

